/*
 * Copyright 2020 Google LLC
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *      http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

`DEFINE_FC_INSTR(C_FLD, CL_FORMAT, LOAD, RV32DC, UIMM)
`DEFINE_FC_INSTR(C_FSD, CS_FORMAT, STORE, RV32DC, UIMM)
`DEFINE_FC_INSTR(C_FLDSP, CI_FORMAT, LOAD, RV32DC, UIMM)
`DEFINE_FC_INSTR(C_FSDSP, CSS_FORMAT, STORE, RV32DC, UIMM)
