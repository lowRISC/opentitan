../../top_earlgrey/rtl/usr_access_xil7series.sv