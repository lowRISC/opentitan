// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "rstmgr_base_vseq.sv"
`include "rstmgr_por_stretcher_vseq.sv"
`include "rstmgr_reset_vseq.sv"
`include "rstmgr_smoke_vseq.sv"
`include "rstmgr_stress_all_vseq.sv"
`include "rstmgr_sw_rst_reset_race_vseq.sv"
`include "rstmgr_sw_rst_vseq.sv"
`include "rstmgr_common_vseq.sv"
`include "rstmgr_sec_cm_scan_intersig_mubi_vseq.sv"
`include "rstmgr_leaf_rst_cnsty_vseq.sv"
`include "rstmgr_leaf_rst_shadow_attack_vseq.sv"
