// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

// Basic sanity test

class ibex_icache_sanity_vseq extends ibex_icache_base_vseq;

  `uvm_object_utils(ibex_icache_sanity_vseq)
  `uvm_object_new

  // No customisation of base class needed

endclass : ibex_icache_sanity_vseq
