// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "flash_ctrl_base_vseq.sv"
`include "flash_ctrl_common_vseq.sv"
`include "flash_ctrl_rand_ops_vseq.sv"
`include "flash_ctrl_smoke_vseq.sv"
