`DEFINE_FP_INSTR(FCVT_L_S,  I_FORMAT, ARITHMETIC, RV64F)
`DEFINE_FP_INSTR(FCVT_LU_S, I_FORMAT, ARITHMETIC, RV64F)
`DEFINE_FP_INSTR(FCVT_S_L,  I_FORMAT, ARITHMETIC, RV64F)
`DEFINE_FP_INSTR(FCVT_S_LU, I_FORMAT, ARITHMETIC, RV64F)
