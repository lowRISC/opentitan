// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "alert_handler_base_vseq.sv"
`include "alert_handler_smoke_vseq.sv"
`include "alert_handler_common_vseq.sv"
`include "alert_handler_random_alerts_vseq.sv"
`include "alert_handler_random_classes_vseq.sv"
`include "alert_handler_esc_intr_timeout_vseq.sv"
`include "alert_handler_esc_alert_accum_vseq.sv"
`include "alert_handler_sig_int_fail_vseq.sv"
`include "alert_handler_entropy_vseq.sv"
`include "alert_handler_ping_timeout_vseq.sv"
`include "alert_handler_lpg_vseq.sv"
`include "alert_handler_lpg_stub_clk_vseq.sv"
`include "alert_handler_stress_all_vseq.sv"
