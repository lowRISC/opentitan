// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "sysrst_ctrl_base_seq.sv"
`include "sysrst_ctrl_in_out_passthrough_seq.sv"

