// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "jtag_riscv_base_seq.sv"
`include "jtag_riscv_csr_seq.sv"
`include "jtag_riscv_dm_activation_seq.sv"
