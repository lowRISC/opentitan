// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "push_pull_base_seq.sv"
`include "push_pull_host_seq.sv"
`include "push_pull_device_seq.sv"
