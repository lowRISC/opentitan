// Copyright lowRISC contributors (OpenTitan project).
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "otp_ctrl_callback_vseq.sv"
`include "otp_ctrl_base_vseq.sv"
`include "otp_ctrl_wake_up_vseq.sv"
`include "otp_ctrl_smoke_vseq.sv"
`include "otp_ctrl_common_vseq.sv"
`include "otp_ctrl_partition_walk_vseq.sv"
`include "otp_ctrl_low_freq_read_vseq.sv"
`include "otp_ctrl_init_fail_vseq.sv"
`include "otp_ctrl_dai_lock_vseq.sv"
`include "otp_ctrl_dai_errs_vseq.sv"
`include "otp_ctrl_macro_errs_vseq.sv"
`include "otp_ctrl_background_chks_vseq.sv"
`include "otp_ctrl_check_fail_vseq.sv"
`include "otp_ctrl_parallel_base_vseq.sv"
`include "otp_ctrl_parallel_key_req_vseq.sv"
`include "otp_ctrl_parallel_lc_req_vseq.sv"
`include "otp_ctrl_parallel_lc_esc_vseq.sv"
`include "otp_ctrl_regwen_vseq.sv"
`include "otp_ctrl_test_access_vseq.sv"
`include "otp_ctrl_stress_all_vseq.sv"
