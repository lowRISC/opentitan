`DEFINE_FC_INSTR(C_FLW,   CL_FORMAT, LOAD, RV32FC, UIMM)
`DEFINE_FC_INSTR(C_FSW,   CS_FORMAT, STORE, RV32FC, UIMM)
`DEFINE_FC_INSTR(C_FLWSP, CI_FORMAT, LOAD, RV32FC, UIMM)
`DEFINE_FC_INSTR(C_FSWSP, CSS_FORMAT, STORE, RV32FC, UIMM)
