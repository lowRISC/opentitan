// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "ibex_icache_base_vseq.sv"
`include "ibex_icache_sanity_vseq.sv"
`include "ibex_icache_passthru_vseq.sv"
`include "ibex_icache_caching_vseq.sv"
`include "ibex_icache_invalidation_vseq.sv"
`include "ibex_icache_oldval_vseq.sv"
`include "ibex_icache_back_line_vseq.sv"
`include "ibex_icache_many_errors_vseq.sv"
