// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "uart_base_seq.sv"
`include "uart_seq.sv"
`include "uart_default_seq.sv"
