// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

class chip_sw_usbdev_suspend_vseq extends chip_sw_usbdev_dpi_vseq;
  `uvm_object_utils(chip_sw_usbdev_suspend_vseq)

  `uvm_object_new

  virtual task body();
    super.body();
  endtask

endclass : chip_sw_usbdev_suspend_vseq
