// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

class ibex_icache_item extends uvm_sequence_item;

  // random variables

  `uvm_object_utils_begin(ibex_icache_item)
  `uvm_object_utils_end

  `uvm_object_new

endclass
