// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "chip_base_vseq.sv"
`include "chip_common_vseq.sv"
`include "chip_sw_base_vseq.sv"
`include "chip_sw_uart_tx_rx_vseq.sv"
`include "chip_sw_gpio_vseq.sv"
