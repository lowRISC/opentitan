// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

// customized tl seq for CIP
`include "cip_tl_seq_item.sv"

// vseqs
`include "cip_base_vseq.sv"
