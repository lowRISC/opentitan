// TODO: Add custom instruction name enum
CUSTOM_1,
