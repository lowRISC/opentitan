`DEFINE_C_INSTR(C_SRLI64, CB_FORMAT, SHIFT, RV128C, NZUIMM)
`DEFINE_C_INSTR(C_SRAI64, CB_FORMAT, SHIFT, RV128C, NZUIMM)
`DEFINE_C_INSTR(C_SLLI64, CI_FORMAT, SHIFT, RV128C, NZUIMM)
`DEFINE_C_INSTR(C_LQ,     CL_FORMAT, LOAD, RV32DC, UIMM)
`DEFINE_C_INSTR(C_SQ,     CS_FORMAT, STORE, RV32DC, UIMM)
`DEFINE_C_INSTR(C_LQSP,   CI_FORMAT, LOAD, RV32DC, UIMM)
`DEFINE_C_INSTR(C_SQSP,   CSS_FORMAT, STORE, RV32DC, UIMM)
