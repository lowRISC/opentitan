// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "kmac_app_base_seq.sv"
`include "kmac_app_host_seq.sv"
`include "kmac_app_device_seq.sv"
