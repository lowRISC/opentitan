../../top_earlgrey/rtl/clkgen_xil7series.sv