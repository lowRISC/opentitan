`DEFINE_C_INSTR(C_ADDIW,  CI_FORMAT, ARITHMETIC, RV64C)
`DEFINE_C_INSTR(C_SUBW,   CA_FORMAT, ARITHMETIC, RV64C)
`DEFINE_C_INSTR(C_ADDW,   CA_FORMAT, ARITHMETIC, RV64C)
`DEFINE_C_INSTR(C_LD,     CL_FORMAT, LOAD, RV64C, UIMM)
`DEFINE_C_INSTR(C_SD,     CS_FORMAT, STORE, RV64C, UIMM)
`DEFINE_C_INSTR(C_LDSP,   CI_FORMAT, LOAD, RV64C, UIMM)
`DEFINE_C_INSTR(C_SDSP,   CSS_FORMAT, STORE, RV64C, UIMM)
