../../top_earlgrey/rtl/physical_pads.sv