`DEFINE_AMO_INSTR(LR_W,      R_FORMAT, LOAD, RV32A)
`DEFINE_AMO_INSTR(SC_W,      R_FORMAT, STORE, RV32A)
`DEFINE_AMO_INSTR(AMOSWAP_W, R_FORMAT, AMO, RV32A)
`DEFINE_AMO_INSTR(AMOADD_W,  R_FORMAT, AMO, RV32A)
`DEFINE_AMO_INSTR(AMOAND_W,  R_FORMAT, AMO, RV32A)
`DEFINE_AMO_INSTR(AMOOR_W,   R_FORMAT, AMO, RV32A)
`DEFINE_AMO_INSTR(AMOXOR_W,  R_FORMAT, AMO, RV32A)
`DEFINE_AMO_INSTR(AMOMIN_W,  R_FORMAT, AMO, RV32A)
`DEFINE_AMO_INSTR(AMOMAX_W,  R_FORMAT, AMO, RV32A)
`DEFINE_AMO_INSTR(AMOMINU_W, R_FORMAT, AMO, RV32A)
`DEFINE_AMO_INSTR(AMOMAXU_W, R_FORMAT, AMO, RV32A)
