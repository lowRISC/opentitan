`include "ibex_asm_program_gen.sv"
`include "ibex_directed_instr_lib.sv"
`include "ibex_debug_triggers_overrides.sv"
