// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`ifndef DATE_DPI_SVH
`define DATE_DPI_SVH

import "DPI-C" function longint get_unix_timestamp();

`endif
