// Copyright lowRISC contributors (OpenTitan project).
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "ac_range_check_base_vseq.sv"
`include "ac_range_check_smoke_vseq.sv"
`include "ac_range_check_smoke_racl_vseq.sv"
`include "ac_range_check_bypass_vseq.sv"
`include "ac_range_check_lock_range_vseq.sv"
`include "ac_range_check_common_vseq.sv"
`include "ac_range_check_stress_all_vseq.sv"
