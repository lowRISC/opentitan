`DEFINE_FP_INSTR(FMV_X_D,   I_FORMAT, ARITHMETIC, RV64D)
`DEFINE_FP_INSTR(FMV_D_X,   I_FORMAT, ARITHMETIC, RV64D)
`DEFINE_FP_INSTR(FCVT_L_D,  I_FORMAT, ARITHMETIC, RV64D)
`DEFINE_FP_INSTR(FCVT_LU_D, I_FORMAT, ARITHMETIC, RV64D)
`DEFINE_FP_INSTR(FCVT_D_L,  I_FORMAT, ARITHMETIC, RV64D)
`DEFINE_FP_INSTR(FCVT_D_LU, I_FORMAT, ARITHMETIC, RV64D)
