`DEFINE_FC_INSTR(C_FLD,   CL_FORMAT, LOAD, RV32DC, UIMM)
`DEFINE_FC_INSTR(C_FSD,   CS_FORMAT, STORE, RV32DC, UIMM)
`DEFINE_FC_INSTR(C_FLDSP, CI_FORMAT, LOAD, RV32DC, UIMM)
`DEFINE_FC_INSTR(C_FSDSP, CSS_FORMAT, STORE, RV32DC, UIMM)
