// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

class spi_sequencer extends dv_seq_sequencer#(spi_item, spi_agent_cfg);
  `uvm_component_utils(spi_sequencer)

  `uvm_component_new

endclass : spi_sequencer
