////////////  RV32M instructions  //////////////
`DEFINE_INSTR(MUL,    R_FORMAT, ARITHMETIC, RV32M)
`DEFINE_INSTR(MULH,   R_FORMAT, ARITHMETIC, RV32M)
`DEFINE_INSTR(MULHSU, R_FORMAT, ARITHMETIC, RV32M)
`DEFINE_INSTR(MULHU,  R_FORMAT, ARITHMETIC, RV32M)
`DEFINE_INSTR(DIV,    R_FORMAT, ARITHMETIC, RV32M)
`DEFINE_INSTR(DIVU,   R_FORMAT, ARITHMETIC, RV32M)
`DEFINE_INSTR(REM,    R_FORMAT, ARITHMETIC, RV32M)
`DEFINE_INSTR(REMU,   R_FORMAT, ARITHMETIC, RV32M)
