../../top_earlgrey/rtl/padring.sv