// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

interface usb20_if ();

  // interface pins
  logic dp;
  logic dm;
  logic tx_mode;
  logic vbus;
  logic susp;
  logic dp_pullup;
  logic dm_pullup;

  // debug signals

endinterface
