// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

class alert_sequencer extends dv_base_sequencer#(alert_seq_item, alert_agent_cfg);
  `uvm_component_utils(alert_sequencer)

  `uvm_component_new

endclass
