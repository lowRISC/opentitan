// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

package alert_handler_test_pkg;
  // dep packages
  import uvm_pkg::*;
  import cip_base_pkg::*;
  import alert_handler_env_pkg::*;

  // macro includes
  `include "uvm_macros.svh"
  `include "dv_macros.svh"

  // local types

  // functions

  // package sources
  `include "alert_handler_base_test.sv"

endpackage
