// Copyright lowRISC contributors (OpenTitan project).
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
package chip_test_pkg;
  // dep packages
  import uvm_pkg::*;
  import cip_base_pkg::*;
  import chip_common_pkg::*;
  import chip_env_pkg::*;
  import tl_agent_pkg::*;

  // macro includes
  `include "uvm_macros.svh"
  `include "dv_macros.svh"

  // local types

  // functions

  // package sources
  `include "chip_base_test.sv"

endpackage
