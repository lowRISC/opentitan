// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

localparam int unsigned DATA_IND_OP_COUNT = 'd37;
