// Copyright lowRISC contributors (OpenTitan project).
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

package top_pkg;

localparam int TL_AW=32;
localparam int TL_DW=32;    // = TL_DBW * 8; TL_DBW must be a power-of-two
localparam int TL_AIW=8;    // a_source, d_source
localparam int TL_DIW=1;    // d_sink
localparam int TL_AUW=21;   // a_user
localparam int TL_DUW=14;   // d_user
localparam int TL_DBW=(TL_DW>>3);
localparam int TL_SZW=$clog2($clog2(TL_DBW)+1);

// Datapath width from the entropy source IP to the actual source of randomness.
// This parameter is top-specific and depends on the actully used source of randomness.
parameter int RNG_BUS_WIDTH = 16;

// NOTE THAT THIS IS A FEATURE FOR TEST CHIPS ONLY TO MITIGATE
// THE RISK OF A BROKEN OTP MACRO. THIS WILL BE DISABLED FOR
// PRODUCTION DEVICES.
localparam int SecVolatileRawUnlockEn = 1;

// The CTN SRAM is set to the same size as the discrete flash (2 x 512kB).
localparam int CtnSramSize = 2 * 512 * 1024;
localparam int CtnSramDepth = CtnSramSize / TL_DBW;
localparam int CtnSramAw = prim_util_pkg::vbits(CtnSramDepth);

endpackage
