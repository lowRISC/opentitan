// Copyright lowRISC contributors (OpenTitan project).
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

class csrng_host_driver extends csrng_driver;
  `uvm_component_utils(csrng_host_driver)
  `uvm_component_new

  // Break down the data and send it to push_pull_host_driver through its sequencer
  csrng_sequencer   m_csrng_sequencer;

  // reset signals
  virtual task reset_signals();
//    `uvm_fatal(`gtn, "FIXME")
  endtask

  // drive trans received from sequencer
  virtual task get_and_drive();
    forever begin
      seq_item_port.get_next_item(req);
      $cast(rsp, req.clone());
      rsp.set_id_info(req);
      `uvm_info(`gfn, $sformatf("rcvd item:\n%0s", req.sprint()), UVM_HIGH)
      // TODO: do the driving part
      //
      // send rsp back to seq
      `uvm_info(`gfn, "item sent", UVM_HIGH)
      seq_item_port.item_done(rsp);
    end
  endtask

endclass
