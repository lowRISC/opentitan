// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "i2c_base_seq.sv"
`include "i2c_device_response_seq.sv"
`include "i2c_target_base_seq.sv"
`include "i2c_target_may_nack_seq.sv"
