// Add your custom extensions, you can list all your local extended SV files here
