// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "key_sideload_base_seq.sv"
`include "key_sideload_set_seq.sv"
