// Copyright lowRISC contributors (OpenTitan project).
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

class chip_sw_ast_clk_outputs_vseq extends chip_sw_base_vseq;
  `uvm_object_utils(chip_sw_ast_clk_outputs_vseq)

  `uvm_object_new

  task body();
     super.body();
  endtask // body

endclass
