`include "ibex_asm_program_gen.sv"
