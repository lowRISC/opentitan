`DEFINE_AMO_INSTR(LR_D,      R_FORMAT, LOAD, RV64A)
`DEFINE_AMO_INSTR(SC_D,      R_FORMAT, STORE, RV64A)
`DEFINE_AMO_INSTR(AMOSWAP_D, R_FORMAT, AMO, RV64A)
`DEFINE_AMO_INSTR(AMOADD_D,  R_FORMAT, AMO, RV64A)
`DEFINE_AMO_INSTR(AMOAND_D,  R_FORMAT, AMO, RV64A)
`DEFINE_AMO_INSTR(AMOOR_D,   R_FORMAT, AMO, RV64A)
`DEFINE_AMO_INSTR(AMOXOR_D,  R_FORMAT, AMO, RV64A)
`DEFINE_AMO_INSTR(AMOMIN_D,  R_FORMAT, AMO, RV64A)
`DEFINE_AMO_INSTR(AMOMAX_D,  R_FORMAT, AMO, RV64A)
`DEFINE_AMO_INSTR(AMOMINU_D, R_FORMAT, AMO, RV64A)
`DEFINE_AMO_INSTR(AMOMAXU_D, R_FORMAT, AMO, RV64A)
