// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "tl_host_base_seq.sv"
`include "tl_host_seq.sv"
`include "tl_host_single_seq.sv"
`include "tl_host_custom_seq.sv"
`include "tl_host_protocol_err_seq.sv"
`include "tl_device_seq.sv"
