// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
// Pseudo driver to access CSR via JTAG TAP
class jtag_riscv_driver extends dv_base_driver #(jtag_riscv_item, jtag_riscv_agent_cfg);

  // drive_jtag process handle
  protected process m_drive_jtag_process_h;

  `uvm_object_utils(jtag_riscv_driver)

  `uvm_object_new

  // reset signals
  virtual task reset_signals();
    `uvm_info(`gfn, "reset_signals: STARTED", UVM_MEDIUM)
    // Kill drive_jtag if its running
    if(m_drive_jtag_process_h != null) m_drive_jtag_process_h.kill();
    // Kill any sequences running on the physical jtag sequencer
    cfg.jtag_sequencer_h.stop_sequences();
  endtask

  // drive trans received from sequencer
  protected virtual task get_and_drive();
    `uvm_info(`gfn, "get_and_drive: STARTED", UVM_MEDIUM)
    forever begin
      seq_item_port.get_next_item(req);
      `uvm_info(`gfn, {"got request: ", req.sprint(uvm_default_line_printer)}, UVM_HIGH)
      accept_tr(req);
      `downcast(rsp, req.clone())
      rsp.set_id_info(req);
      seq_item_port.item_done();
      fork
        begin : drive_jtag_process
          m_drive_jtag_process_h = process::self();
          drive_jtag(rsp);
        end : drive_jtag_process
      join
      // Send response
      seq_item_port.put_response(rsp);
    end
  endtask

  protected virtual task drive_jtag(ITEM_T drive_req);
    bit [DMI_DATAW-1:0] dout;
    bit [DMI_DATAW-1:0] rdata;
    bit [DMI_OPW-1:0] status;

    `uvm_info(`gfn, {"drive_jtag: ",
         drive_req.sprint(uvm_default_line_printer)}, UVM_HIGH)

    // Mark start of transaction processing
    void'(begin_tr(drive_req));

    // Drive IR with DMI access
    send_riscv_ir_req(JtagDmiAccess);

    // Drive DR with operation type, address, and data
    send_csr_dr_req(drive_req.op, drive_req.data, drive_req.addr, dout);

    // Get status of previous transfer
    check_csr_req_status(status, rdata);
    drive_req.status = status;

    // Update CSR read data
    if (drive_req.op == DmiRead) drive_req.data = rdata;

    // Mark end of transaction processing
    end_tr(drive_req);

  endtask

 protected virtual task send_riscv_ir_req(jtag_ir_e riscv_ir_req);
    jtag_ir_seq ir_seq;
    `uvm_create_obj(jtag_ir_seq, ir_seq);
    `DV_CHECK_RANDOMIZE_WITH_FATAL(ir_seq,
        ir_len == DMI_IRW;
        ir     == riscv_ir_req;)
    ir_seq.start(cfg.jtag_sequencer_h);
  endtask

  protected virtual task send_dtmcs_dr_req(jtag_dtmcs_e dtmcs_req_idx);
    jtag_dr_seq dr_seq;
    `uvm_create_obj(jtag_dr_seq, dr_seq);
    `DV_CHECK_RANDOMIZE_WITH_FATAL(dr_seq,
        dr_len == DTMCS_DRW;
        dr     == 1 << dtmcs_req_idx;)
    dr_seq.start(cfg.jtag_sequencer_h);
  endtask

  // This task sends a CSR register read/write request via JTAG data register.
  protected virtual task send_csr_dr_req(input bit [DMI_OPW-1:0]    op,
                               input bit [DMI_DATAW-1:0]  data,
                               input bit [DMI_ADDRW-1:0]  addr,
                               output bit [DMI_DATAW-1:0] dout);
    jtag_dr_seq dr_seq;
    `uvm_create_obj(jtag_dr_seq, dr_seq);
    `DV_CHECK_RANDOMIZE_WITH_FATAL(dr_seq,
        dr_len == DMI_DRW;
        dr     == {addr, data, op};)
    dr_seq.start(cfg.jtag_sequencer_h);
    dout = dr_seq.rsp.dout;
  endtask

  // This task checks a CSR register read/write request status via data request.
  // This task will output operation status and rdata (this rdata is only meaningful if it is a
  // read operation).
  protected virtual task check_csr_req_status(
      ref bit [DMI_OPW-1:0] status, ref bit [DMI_DATAW-1:0] rdata);
    while (1) begin
      bit [DMI_DRW-1:0] dout;
      send_csr_dr_req(DmiStatus, 0, 0, dout);
      status = dout[0 +: DMI_OPW];

      // The DmiInProgress status is sticky and has to be cleared by dmireset via DTMCS.
      if (status == DmiInProgress) begin
        send_riscv_ir_req(JtagDtmCsr);
        send_dtmcs_dr_req(DmiReset);
        send_riscv_ir_req(JtagDmiAccess);
      end

      if (status != DmiInProgress) begin
        rdata = dout[2 +: DMI_DATAW];
        break;
      end
    end
  endtask
endclass
