../../top_earlgrey/rtl/top_pkg.sv