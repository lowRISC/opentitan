// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "keymgr_kmac_base_seq.sv"
`include "keymgr_kmac_host_seq.sv"
`include "keymgr_kmac_device_seq.sv"
