class usb20_sequencer extends dv_base_sequencer#( usb20_item, usb20_agent_cfg);
  
    `uvm_sequencer_utils(usb20_sequencer)
    `uvm_component_new 
    
endclass : usb20_sequencer
