// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "spi_base_seq.sv"
`include "spi_host_seq.sv"
`include "spi_host_flash_seq.sv"
`include "spi_host_tpm_seq.sv"
`include "spi_device_flash_seq.sv"
`include "spi_host_dummy_seq.sv"
`include "spi_device_seq.sv"
`include "spi_device_cmd_rsp_seq.sv"
