// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

class csrng_item extends uvm_sequence_item;

  // TODO: create
  `uvm_object_utils_begin(csrng_item)
  `uvm_object_utils_end

  `uvm_object_new

endclass
