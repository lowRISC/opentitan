`DEFINE_INSTR(MULW,   R_FORMAT, ARITHMETIC, RV64M)
`DEFINE_INSTR(DIVW,   R_FORMAT, ARITHMETIC, RV64M)
`DEFINE_INSTR(DIVUW,  R_FORMAT, ARITHMETIC, RV64M)
`DEFINE_INSTR(REMW,   R_FORMAT, ARITHMETIC, RV64M)
`DEFINE_INSTR(REMUW,  R_FORMAT, ARITHMETIC, RV64M)
